-- Computer_System_VGA_Subsystem_Char_Buf_Subsystem.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Computer_System_VGA_Subsystem_Char_Buf_Subsystem is
	port (
		avalon_char_source_ready             : in  std_logic                     := '0';             --        avalon_char_source.ready
		avalon_char_source_startofpacket     : out std_logic;                                        --                          .startofpacket
		avalon_char_source_endofpacket       : out std_logic;                                        --                          .endofpacket
		avalon_char_source_valid             : out std_logic;                                        --                          .valid
		avalon_char_source_data              : out std_logic_vector(39 downto 0);                    --                          .data
		char_buffer_control_slave_address    : in  std_logic_vector(1 downto 0)  := (others => '0'); -- char_buffer_control_slave.address
		char_buffer_control_slave_byteenable : in  std_logic_vector(3 downto 0)  := (others => '0'); --                          .byteenable
		char_buffer_control_slave_read       : in  std_logic                     := '0';             --                          .read
		char_buffer_control_slave_write      : in  std_logic                     := '0';             --                          .write
		char_buffer_control_slave_writedata  : in  std_logic_vector(31 downto 0) := (others => '0'); --                          .writedata
		char_buffer_control_slave_readdata   : out std_logic_vector(31 downto 0);                    --                          .readdata
		char_buffer_slave_address            : in  std_logic_vector(10 downto 0) := (others => '0'); --         char_buffer_slave.address
		char_buffer_slave_clken              : in  std_logic                     := '0';             --                          .clken
		char_buffer_slave_chipselect         : in  std_logic                     := '0';             --                          .chipselect
		char_buffer_slave_write              : in  std_logic                     := '0';             --                          .write
		char_buffer_slave_readdata           : out std_logic_vector(31 downto 0);                    --                          .readdata
		char_buffer_slave_writedata          : in  std_logic_vector(31 downto 0) := (others => '0'); --                          .writedata
		char_buffer_slave_byteenable         : in  std_logic_vector(3 downto 0)  := (others => '0'); --                          .byteenable
		sys_clk_clk                          : in  std_logic                     := '0';             --                   sys_clk.clk
		sys_reset_reset_n                    : in  std_logic                     := '0'              --                 sys_reset.reset_n
	);
end entity Computer_System_VGA_Subsystem_Char_Buf_Subsystem;

architecture rtl of Computer_System_VGA_Subsystem_Char_Buf_Subsystem is
	component Computer_System_VGA_Subsystem_Char_Buf_Subsystem_ASCII_to_Image is
		port (
			clk                     : in  std_logic                    := 'X';             -- clk
			reset                   : in  std_logic                    := 'X';             -- reset
			ascii_in_channel        : in  std_logic_vector(5 downto 0) := (others => 'X'); -- channel
			ascii_in_startofpacket  : in  std_logic                    := 'X';             -- startofpacket
			ascii_in_endofpacket    : in  std_logic                    := 'X';             -- endofpacket
			ascii_in_valid          : in  std_logic                    := 'X';             -- valid
			ascii_in_ready          : out std_logic;                                       -- ready
			ascii_in_data           : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			image_out_ready         : in  std_logic                    := 'X';             -- ready
			image_out_startofpacket : out std_logic;                                       -- startofpacket
			image_out_endofpacket   : out std_logic;                                       -- endofpacket
			image_out_valid         : out std_logic;                                       -- valid
			image_out_data          : out std_logic                                        -- data
		);
	end component Computer_System_VGA_Subsystem_Char_Buf_Subsystem_ASCII_to_Image;

	component Computer_System_VGA_Subsystem_Char_Buf_Subsystem_Char_Buf_DMA is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_arbiterlock   : out std_logic;                                        -- lock
			master_read          : out std_logic;                                        -- read
			master_readdata      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_data          : out std_logic_vector(7 downto 0);                     -- data
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic                                         -- valid
		);
	end component Computer_System_VGA_Subsystem_Char_Buf_Subsystem_Char_Buf_DMA;

	component Computer_System_VGA_Subsystem_Char_Buf_Subsystem_Char_Buf_RGB_Resampler is
		port (
			clk                      : in  std_logic                     := 'X'; -- clk
			reset                    : in  std_logic                     := 'X'; -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X'; -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X'; -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X'; -- valid
			stream_in_ready          : out std_logic;                            -- ready
			stream_in_data           : in  std_logic                     := 'X'; -- data
			slave_read               : in  std_logic                     := 'X'; -- read
			slave_readdata           : out std_logic_vector(31 downto 0);        -- readdata
			stream_out_ready         : in  std_logic                     := 'X'; -- ready
			stream_out_startofpacket : out std_logic;                            -- startofpacket
			stream_out_endofpacket   : out std_logic;                            -- endofpacket
			stream_out_valid         : out std_logic;                            -- valid
			stream_out_data          : out std_logic_vector(39 downto 0)         -- data
		);
	end component Computer_System_VGA_Subsystem_Char_Buf_Subsystem_Char_Buf_RGB_Resampler;

	component Computer_System_VGA_Subsystem_Char_Buf_Subsystem_Char_Buf_Scaler is
		port (
			clk                      : in  std_logic                    := 'X';             -- clk
			reset                    : in  std_logic                    := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                    := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                    := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                    := 'X';             -- valid
			stream_in_ready          : out std_logic;                                       -- ready
			stream_in_data           : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                    := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                       -- startofpacket
			stream_out_endofpacket   : out std_logic;                                       -- endofpacket
			stream_out_valid         : out std_logic;                                       -- valid
			stream_out_data          : out std_logic_vector(7 downto 0);                    -- data
			stream_out_channel       : out std_logic_vector(5 downto 0)                     -- channel
		);
	end component Computer_System_VGA_Subsystem_Char_Buf_Subsystem_Char_Buf_Scaler;

	component Computer_System_VGA_Subsystem_Char_Buf_Subsystem_Onchip_SRAM is
		port (
			address     : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			address2    : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk         : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			freeze      : in  std_logic                     := 'X'              -- freeze
		);
	end component Computer_System_VGA_Subsystem_Char_Buf_Subsystem_Onchip_SRAM;

	component Computer_System_VGA_Subsystem_Char_Buf_Subsystem_Set_Black_Transparent is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(39 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(39 downto 0)                     -- data
		);
	end component Computer_System_VGA_Subsystem_Char_Buf_Subsystem_Set_Black_Transparent;

	component Computer_System_VGA_Subsystem_Char_Buf_Subsystem_mm_interconnect_0 is
		port (
			Sys_Clk_clk_clk                                : in  std_logic                     := 'X';             -- clk
			Char_Buf_DMA_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			Char_Buf_DMA_avalon_dma_master_address         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			Char_Buf_DMA_avalon_dma_master_waitrequest     : out std_logic;                                        -- waitrequest
			Char_Buf_DMA_avalon_dma_master_read            : in  std_logic                     := 'X';             -- read
			Char_Buf_DMA_avalon_dma_master_readdata        : out std_logic_vector(7 downto 0);                     -- readdata
			Char_Buf_DMA_avalon_dma_master_readdatavalid   : out std_logic;                                        -- readdatavalid
			Char_Buf_DMA_avalon_dma_master_lock            : in  std_logic                     := 'X';             -- lock
			Onchip_SRAM_s2_address                         : out std_logic_vector(10 downto 0);                    -- address
			Onchip_SRAM_s2_write                           : out std_logic;                                        -- write
			Onchip_SRAM_s2_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Onchip_SRAM_s2_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			Onchip_SRAM_s2_byteenable                      : out std_logic_vector(3 downto 0);                     -- byteenable
			Onchip_SRAM_s2_chipselect                      : out std_logic;                                        -- chipselect
			Onchip_SRAM_s2_clken                           : out std_logic                                         -- clken
		);
	end component Computer_System_VGA_Subsystem_Char_Buf_Subsystem_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal ascii_to_image_avalon_image_source_valid               : std_logic;                     -- ASCII_to_Image:image_out_valid -> Char_Buf_RGB_Resampler:stream_in_valid
	signal ascii_to_image_avalon_image_source_data                : std_logic;                     -- ASCII_to_Image:image_out_data -> Char_Buf_RGB_Resampler:stream_in_data
	signal ascii_to_image_avalon_image_source_ready               : std_logic;                     -- Char_Buf_RGB_Resampler:stream_in_ready -> ASCII_to_Image:image_out_ready
	signal ascii_to_image_avalon_image_source_startofpacket       : std_logic;                     -- ASCII_to_Image:image_out_startofpacket -> Char_Buf_RGB_Resampler:stream_in_startofpacket
	signal ascii_to_image_avalon_image_source_endofpacket         : std_logic;                     -- ASCII_to_Image:image_out_endofpacket -> Char_Buf_RGB_Resampler:stream_in_endofpacket
	signal char_buf_dma_avalon_pixel_source_valid                 : std_logic;                     -- Char_Buf_DMA:stream_valid -> Char_Buf_Scaler:stream_in_valid
	signal char_buf_dma_avalon_pixel_source_data                  : std_logic_vector(7 downto 0);  -- Char_Buf_DMA:stream_data -> Char_Buf_Scaler:stream_in_data
	signal char_buf_dma_avalon_pixel_source_ready                 : std_logic;                     -- Char_Buf_Scaler:stream_in_ready -> Char_Buf_DMA:stream_ready
	signal char_buf_dma_avalon_pixel_source_startofpacket         : std_logic;                     -- Char_Buf_DMA:stream_startofpacket -> Char_Buf_Scaler:stream_in_startofpacket
	signal char_buf_dma_avalon_pixel_source_endofpacket           : std_logic;                     -- Char_Buf_DMA:stream_endofpacket -> Char_Buf_Scaler:stream_in_endofpacket
	signal char_buf_rgb_resampler_avalon_rgb_source_valid         : std_logic;                     -- Char_Buf_RGB_Resampler:stream_out_valid -> Set_Black_Transparent:stream_in_valid
	signal char_buf_rgb_resampler_avalon_rgb_source_data          : std_logic_vector(39 downto 0); -- Char_Buf_RGB_Resampler:stream_out_data -> Set_Black_Transparent:stream_in_data
	signal char_buf_rgb_resampler_avalon_rgb_source_ready         : std_logic;                     -- Set_Black_Transparent:stream_in_ready -> Char_Buf_RGB_Resampler:stream_out_ready
	signal char_buf_rgb_resampler_avalon_rgb_source_startofpacket : std_logic;                     -- Char_Buf_RGB_Resampler:stream_out_startofpacket -> Set_Black_Transparent:stream_in_startofpacket
	signal char_buf_rgb_resampler_avalon_rgb_source_endofpacket   : std_logic;                     -- Char_Buf_RGB_Resampler:stream_out_endofpacket -> Set_Black_Transparent:stream_in_endofpacket
	signal char_buf_scaler_avalon_scaler_source_valid             : std_logic;                     -- Char_Buf_Scaler:stream_out_valid -> ASCII_to_Image:ascii_in_valid
	signal char_buf_scaler_avalon_scaler_source_data              : std_logic_vector(7 downto 0);  -- Char_Buf_Scaler:stream_out_data -> ASCII_to_Image:ascii_in_data
	signal char_buf_scaler_avalon_scaler_source_ready             : std_logic;                     -- ASCII_to_Image:ascii_in_ready -> Char_Buf_Scaler:stream_out_ready
	signal char_buf_scaler_avalon_scaler_source_channel           : std_logic_vector(5 downto 0);  -- Char_Buf_Scaler:stream_out_channel -> ASCII_to_Image:ascii_in_channel
	signal char_buf_scaler_avalon_scaler_source_startofpacket     : std_logic;                     -- Char_Buf_Scaler:stream_out_startofpacket -> ASCII_to_Image:ascii_in_startofpacket
	signal char_buf_scaler_avalon_scaler_source_endofpacket       : std_logic;                     -- Char_Buf_Scaler:stream_out_endofpacket -> ASCII_to_Image:ascii_in_endofpacket
	signal char_buf_dma_avalon_dma_master_waitrequest             : std_logic;                     -- mm_interconnect_0:Char_Buf_DMA_avalon_dma_master_waitrequest -> Char_Buf_DMA:master_waitrequest
	signal char_buf_dma_avalon_dma_master_readdata                : std_logic_vector(7 downto 0);  -- mm_interconnect_0:Char_Buf_DMA_avalon_dma_master_readdata -> Char_Buf_DMA:master_readdata
	signal char_buf_dma_avalon_dma_master_address                 : std_logic_vector(31 downto 0); -- Char_Buf_DMA:master_address -> mm_interconnect_0:Char_Buf_DMA_avalon_dma_master_address
	signal char_buf_dma_avalon_dma_master_read                    : std_logic;                     -- Char_Buf_DMA:master_read -> mm_interconnect_0:Char_Buf_DMA_avalon_dma_master_read
	signal char_buf_dma_avalon_dma_master_readdatavalid           : std_logic;                     -- mm_interconnect_0:Char_Buf_DMA_avalon_dma_master_readdatavalid -> Char_Buf_DMA:master_readdatavalid
	signal char_buf_dma_avalon_dma_master_lock                    : std_logic;                     -- Char_Buf_DMA:master_arbiterlock -> mm_interconnect_0:Char_Buf_DMA_avalon_dma_master_lock
	signal mm_interconnect_0_onchip_sram_s2_chipselect            : std_logic;                     -- mm_interconnect_0:Onchip_SRAM_s2_chipselect -> Onchip_SRAM:chipselect2
	signal mm_interconnect_0_onchip_sram_s2_readdata              : std_logic_vector(31 downto 0); -- Onchip_SRAM:readdata2 -> mm_interconnect_0:Onchip_SRAM_s2_readdata
	signal mm_interconnect_0_onchip_sram_s2_address               : std_logic_vector(10 downto 0); -- mm_interconnect_0:Onchip_SRAM_s2_address -> Onchip_SRAM:address2
	signal mm_interconnect_0_onchip_sram_s2_byteenable            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:Onchip_SRAM_s2_byteenable -> Onchip_SRAM:byteenable2
	signal mm_interconnect_0_onchip_sram_s2_write                 : std_logic;                     -- mm_interconnect_0:Onchip_SRAM_s2_write -> Onchip_SRAM:write2
	signal mm_interconnect_0_onchip_sram_s2_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:Onchip_SRAM_s2_writedata -> Onchip_SRAM:writedata2
	signal mm_interconnect_0_onchip_sram_s2_clken                 : std_logic;                     -- mm_interconnect_0:Onchip_SRAM_s2_clken -> Onchip_SRAM:clken2
	signal rst_controller_reset_out_reset                         : std_logic;                     -- rst_controller:reset_out -> [ASCII_to_Image:reset, Char_Buf_DMA:reset, Char_Buf_RGB_Resampler:reset, Char_Buf_Scaler:reset, Onchip_SRAM:reset, Set_Black_Transparent:reset, mm_interconnect_0:Char_Buf_DMA_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                     : std_logic;                     -- rst_controller:reset_req -> [Onchip_SRAM:reset_req, rst_translator:reset_req_in]
	signal sys_reset_reset_n_ports_inv                            : std_logic;                     -- sys_reset_reset_n:inv -> rst_controller:reset_in0

begin

	ascii_to_image : component Computer_System_VGA_Subsystem_Char_Buf_Subsystem_ASCII_to_Image
		port map (
			clk                     => sys_clk_clk,                                        --                 clk.clk
			reset                   => rst_controller_reset_out_reset,                     --               reset.reset
			ascii_in_channel        => char_buf_scaler_avalon_scaler_source_channel,       --   avalon_ascii_sink.channel
			ascii_in_startofpacket  => char_buf_scaler_avalon_scaler_source_startofpacket, --                    .startofpacket
			ascii_in_endofpacket    => char_buf_scaler_avalon_scaler_source_endofpacket,   --                    .endofpacket
			ascii_in_valid          => char_buf_scaler_avalon_scaler_source_valid,         --                    .valid
			ascii_in_ready          => char_buf_scaler_avalon_scaler_source_ready,         --                    .ready
			ascii_in_data           => char_buf_scaler_avalon_scaler_source_data,          --                    .data
			image_out_ready         => ascii_to_image_avalon_image_source_ready,           -- avalon_image_source.ready
			image_out_startofpacket => ascii_to_image_avalon_image_source_startofpacket,   --                    .startofpacket
			image_out_endofpacket   => ascii_to_image_avalon_image_source_endofpacket,     --                    .endofpacket
			image_out_valid         => ascii_to_image_avalon_image_source_valid,           --                    .valid
			image_out_data          => ascii_to_image_avalon_image_source_data             --                    .data
		);

	char_buf_dma : component Computer_System_VGA_Subsystem_Char_Buf_Subsystem_Char_Buf_DMA
		port map (
			clk                  => sys_clk_clk,                                    --                      clk.clk
			reset                => rst_controller_reset_out_reset,                 --                    reset.reset
			master_address       => char_buf_dma_avalon_dma_master_address,         --        avalon_dma_master.address
			master_waitrequest   => char_buf_dma_avalon_dma_master_waitrequest,     --                         .waitrequest
			master_arbiterlock   => char_buf_dma_avalon_dma_master_lock,            --                         .lock
			master_read          => char_buf_dma_avalon_dma_master_read,            --                         .read
			master_readdata      => char_buf_dma_avalon_dma_master_readdata,        --                         .readdata
			master_readdatavalid => char_buf_dma_avalon_dma_master_readdatavalid,   --                         .readdatavalid
			slave_address        => char_buffer_control_slave_address,              -- avalon_dma_control_slave.address
			slave_byteenable     => char_buffer_control_slave_byteenable,           --                         .byteenable
			slave_read           => char_buffer_control_slave_read,                 --                         .read
			slave_write          => char_buffer_control_slave_write,                --                         .write
			slave_writedata      => char_buffer_control_slave_writedata,            --                         .writedata
			slave_readdata       => char_buffer_control_slave_readdata,             --                         .readdata
			stream_ready         => char_buf_dma_avalon_pixel_source_ready,         --      avalon_pixel_source.ready
			stream_data          => char_buf_dma_avalon_pixel_source_data,          --                         .data
			stream_startofpacket => char_buf_dma_avalon_pixel_source_startofpacket, --                         .startofpacket
			stream_endofpacket   => char_buf_dma_avalon_pixel_source_endofpacket,   --                         .endofpacket
			stream_valid         => char_buf_dma_avalon_pixel_source_valid          --                         .valid
		);

	char_buf_rgb_resampler : component Computer_System_VGA_Subsystem_Char_Buf_Subsystem_Char_Buf_RGB_Resampler
		port map (
			clk                      => sys_clk_clk,                                            --               clk.clk
			reset                    => rst_controller_reset_out_reset,                         --             reset.reset
			stream_in_startofpacket  => ascii_to_image_avalon_image_source_startofpacket,       --   avalon_rgb_sink.startofpacket
			stream_in_endofpacket    => ascii_to_image_avalon_image_source_endofpacket,         --                  .endofpacket
			stream_in_valid          => ascii_to_image_avalon_image_source_valid,               --                  .valid
			stream_in_ready          => ascii_to_image_avalon_image_source_ready,               --                  .ready
			stream_in_data           => ascii_to_image_avalon_image_source_data,                --                  .data
			slave_read               => open,                                                   --  avalon_rgb_slave.read
			slave_readdata           => open,                                                   --                  .readdata
			stream_out_ready         => char_buf_rgb_resampler_avalon_rgb_source_ready,         -- avalon_rgb_source.ready
			stream_out_startofpacket => char_buf_rgb_resampler_avalon_rgb_source_startofpacket, --                  .startofpacket
			stream_out_endofpacket   => char_buf_rgb_resampler_avalon_rgb_source_endofpacket,   --                  .endofpacket
			stream_out_valid         => char_buf_rgb_resampler_avalon_rgb_source_valid,         --                  .valid
			stream_out_data          => char_buf_rgb_resampler_avalon_rgb_source_data           --                  .data
		);

	char_buf_scaler : component Computer_System_VGA_Subsystem_Char_Buf_Subsystem_Char_Buf_Scaler
		port map (
			clk                      => sys_clk_clk,                                        --                  clk.clk
			reset                    => rst_controller_reset_out_reset,                     --                reset.reset
			stream_in_startofpacket  => char_buf_dma_avalon_pixel_source_startofpacket,     --   avalon_scaler_sink.startofpacket
			stream_in_endofpacket    => char_buf_dma_avalon_pixel_source_endofpacket,       --                     .endofpacket
			stream_in_valid          => char_buf_dma_avalon_pixel_source_valid,             --                     .valid
			stream_in_ready          => char_buf_dma_avalon_pixel_source_ready,             --                     .ready
			stream_in_data           => char_buf_dma_avalon_pixel_source_data,              --                     .data
			stream_out_ready         => char_buf_scaler_avalon_scaler_source_ready,         -- avalon_scaler_source.ready
			stream_out_startofpacket => char_buf_scaler_avalon_scaler_source_startofpacket, --                     .startofpacket
			stream_out_endofpacket   => char_buf_scaler_avalon_scaler_source_endofpacket,   --                     .endofpacket
			stream_out_valid         => char_buf_scaler_avalon_scaler_source_valid,         --                     .valid
			stream_out_data          => char_buf_scaler_avalon_scaler_source_data,          --                     .data
			stream_out_channel       => char_buf_scaler_avalon_scaler_source_channel        --                     .channel
		);

	onchip_sram : component Computer_System_VGA_Subsystem_Char_Buf_Subsystem_Onchip_SRAM
		port map (
			address     => char_buffer_slave_address,                   --     s1.address
			clken       => char_buffer_slave_clken,                     --       .clken
			chipselect  => char_buffer_slave_chipselect,                --       .chipselect
			write       => char_buffer_slave_write,                     --       .write
			readdata    => char_buffer_slave_readdata,                  --       .readdata
			writedata   => char_buffer_slave_writedata,                 --       .writedata
			byteenable  => char_buffer_slave_byteenable,                --       .byteenable
			address2    => mm_interconnect_0_onchip_sram_s2_address,    --     s2.address
			chipselect2 => mm_interconnect_0_onchip_sram_s2_chipselect, --       .chipselect
			clken2      => mm_interconnect_0_onchip_sram_s2_clken,      --       .clken
			write2      => mm_interconnect_0_onchip_sram_s2_write,      --       .write
			readdata2   => mm_interconnect_0_onchip_sram_s2_readdata,   --       .readdata
			writedata2  => mm_interconnect_0_onchip_sram_s2_writedata,  --       .writedata
			byteenable2 => mm_interconnect_0_onchip_sram_s2_byteenable, --       .byteenable
			clk         => sys_clk_clk,                                 --   clk1.clk
			reset       => rst_controller_reset_out_reset,              -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,          --       .reset_req
			freeze      => '0'                                          -- (terminated)
		);

	set_black_transparent : component Computer_System_VGA_Subsystem_Char_Buf_Subsystem_Set_Black_Transparent
		port map (
			clk                      => sys_clk_clk,                                            --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                         --                     reset.reset
			stream_in_startofpacket  => char_buf_rgb_resampler_avalon_rgb_source_startofpacket, --   avalon_apply_alpha_sink.startofpacket
			stream_in_endofpacket    => char_buf_rgb_resampler_avalon_rgb_source_endofpacket,   --                          .endofpacket
			stream_in_valid          => char_buf_rgb_resampler_avalon_rgb_source_valid,         --                          .valid
			stream_in_ready          => char_buf_rgb_resampler_avalon_rgb_source_ready,         --                          .ready
			stream_in_data           => char_buf_rgb_resampler_avalon_rgb_source_data,          --                          .data
			stream_out_ready         => avalon_char_source_ready,                               -- avalon_apply_alpha_source.ready
			stream_out_startofpacket => avalon_char_source_startofpacket,                       --                          .startofpacket
			stream_out_endofpacket   => avalon_char_source_endofpacket,                         --                          .endofpacket
			stream_out_valid         => avalon_char_source_valid,                               --                          .valid
			stream_out_data          => avalon_char_source_data                                 --                          .data
		);

	mm_interconnect_0 : component Computer_System_VGA_Subsystem_Char_Buf_Subsystem_mm_interconnect_0
		port map (
			Sys_Clk_clk_clk                                => sys_clk_clk,                                  --                              Sys_Clk_clk.clk
			Char_Buf_DMA_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,               -- Char_Buf_DMA_reset_reset_bridge_in_reset.reset
			Char_Buf_DMA_avalon_dma_master_address         => char_buf_dma_avalon_dma_master_address,       --           Char_Buf_DMA_avalon_dma_master.address
			Char_Buf_DMA_avalon_dma_master_waitrequest     => char_buf_dma_avalon_dma_master_waitrequest,   --                                         .waitrequest
			Char_Buf_DMA_avalon_dma_master_read            => char_buf_dma_avalon_dma_master_read,          --                                         .read
			Char_Buf_DMA_avalon_dma_master_readdata        => char_buf_dma_avalon_dma_master_readdata,      --                                         .readdata
			Char_Buf_DMA_avalon_dma_master_readdatavalid   => char_buf_dma_avalon_dma_master_readdatavalid, --                                         .readdatavalid
			Char_Buf_DMA_avalon_dma_master_lock            => char_buf_dma_avalon_dma_master_lock,          --                                         .lock
			Onchip_SRAM_s2_address                         => mm_interconnect_0_onchip_sram_s2_address,     --                           Onchip_SRAM_s2.address
			Onchip_SRAM_s2_write                           => mm_interconnect_0_onchip_sram_s2_write,       --                                         .write
			Onchip_SRAM_s2_readdata                        => mm_interconnect_0_onchip_sram_s2_readdata,    --                                         .readdata
			Onchip_SRAM_s2_writedata                       => mm_interconnect_0_onchip_sram_s2_writedata,   --                                         .writedata
			Onchip_SRAM_s2_byteenable                      => mm_interconnect_0_onchip_sram_s2_byteenable,  --                                         .byteenable
			Onchip_SRAM_s2_chipselect                      => mm_interconnect_0_onchip_sram_s2_chipselect,  --                                         .chipselect
			Onchip_SRAM_s2_clken                           => mm_interconnect_0_onchip_sram_s2_clken        --                                         .clken
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => sys_reset_reset_n_ports_inv,        -- reset_in0.reset
			clk            => sys_clk_clk,                        --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	sys_reset_reset_n_ports_inv <= not sys_reset_reset_n;

end architecture rtl; -- of Computer_System_VGA_Subsystem_Char_Buf_Subsystem
